


.SUBCKT sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield

Cx  sky130_fd_pr__cap_vpp_22p5x23p1_pol1m1m2m3m4m5_noshield

.ENDS
