


.SUBCKT sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4 C0 C1 MET4 SUB

Cx C0 C1 MET4 SUB sky130_fd_pr__cap_vpp_06p8x06p1_l1m1m2m3_shieldpom4

.ENDS
