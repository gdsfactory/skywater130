


.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield C0 C1 SUB

Cx C0 C1 SUB sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield

.ENDS
