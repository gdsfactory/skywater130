


.SUBCKT sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3 C0 C1 MET3 SUB

Cx C0 C1 MET3 SUB sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3

.ENDS
