


.SUBCKT sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1 C0 C1 SUB

Cx C0 C1 SUB sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1

.ENDS
