


.SUBCKT sky130_fd_pr__cap_vpp_55p8x23p1_pol1m1m2m3m4m5_noshield_test

Cx  sky130_fd_pr__cap_vpp_55p8x23p1_pol1m1m2m3m4m5_noshield_test

.ENDS
